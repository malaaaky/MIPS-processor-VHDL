`timescale 1ns / 1ps
module datapath(
    input clk, reset,
    input [31:0] instr,
    input [2:0] aluoperation,
    output zero,
    input regwrite,
    input [31:0] aluout
    );


endmodule
